../../../peripheral/src/AddRawFN.sv