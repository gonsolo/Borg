../../../borg_peripheral/src/RoundAnyRawFNToRecFN_ie8_is26_oe8_os24.sv