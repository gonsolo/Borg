../../../borg_peripheral/src/AddRecFN.sv