../../../borg_peripheral/src/RoundRawFNToRecFN_e8_s24.sv