../../../borg_peripheral/src/MulFullRawFN.sv