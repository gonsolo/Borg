../../../borg_peripheral/src/MulAddRecFNToRaw_postMul_e8_s24.sv