../../../peripheral/src/Borg.sv