../../../borg_peripheral/src/MulAddRecFNToRaw_preMul_e8_s24.sv