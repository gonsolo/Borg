../../../borg_peripheral/src/MulRawFN.sv