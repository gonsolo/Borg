../../../borg_peripheral/src/MulRecFN.sv