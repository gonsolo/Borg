../../../borg_peripheral/src/registerFile_4x32.sv