../../../borg_peripheral/src/MulAddRecFN_e8_s24.sv