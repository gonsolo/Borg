../../../borg_peripheral/src/instructionMemory_4x32.sv