../../../borg_peripheral/src/instructionMemory_8x32.sv