../../../borg_peripheral/src/Borg.sv