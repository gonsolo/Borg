../../../borg_peripheral/src/AddRawFN.sv