../../../peripheral/src/AddRecFN.sv